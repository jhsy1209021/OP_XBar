`ifndef XBAR
`define XBAR
    `include "xbar_master_interface.sv"
    `include "xbar_slave_interface.sv"
`endif