`ifndef ASYNC_FIFO_8
`define ASYNC_FIFO_8
    `include "async_fifo_8.sv"
    `include "read_pointer_handler.sv"
    `include "write_pointer_handler.sv"
    `include "graycode_encoder_16.sv"
    `include "synchronizer_3.sv"
`endif