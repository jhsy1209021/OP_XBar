`ifndef ASYNC_FIFO
`define ASYNC_FIFO
    `include "async_fifo.sv"
    `include "read_pointer_handler.sv"
    `include "write_pointer_handler.sv"
    `include "graycode_encoder.sv"
    `include "synchronizer.sv"
`endif