`ifndef XBAR
`define XBAR
    `include "xbar.sv"
    `include "xbar_master_interface.svh"
    `include "xbar_slave_interface.svh"
`endif